library verilog;
use verilog.vl_types.all;
entity spi_test_TB is
end spi_test_TB;
